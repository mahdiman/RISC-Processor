LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE IEEE.math_real.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY writeBack IS
  -- PORT();
END writeBack;

ARCHITECTURE writeBack_arch OF writeBack IS
BEGIN

END writeBack_arch;
